// =============================================================================
// Module  : tb_recurrent_layer
// Description : 재귀 SNN 레이어의 패턴 학습 및 연상 복원 검증
//
// [검증 시나리오]
//
// [학습 단계] 패턴 A = {N0, N1} 동시 발화 반복 학습
//   → W01, W10 강화 기대
//
// [복원 단계] N0만 자극 (패턴의 절반만 입력)
//   → W01이 강화되어 N1도 발화하는지 확인
//   → "N0를 보면 N1이 떠오른다" = 연상 기억!
//
// [관전 포인트]
//   학습 전: N0만 자극 → N0만 발화
//   학습 후: N0만 자극 → N0 + N1 발화 (패턴 복원!)
// =============================================================================
`timescale 1ns / 1ps

module tb_recurrent_layer;

    reg        clk, rst_n;
    reg  [3:0] ext_in;

    wire [3:0] spk;
    wire [7:0] v0, v1, v2, v3;
    wire [7:0] w01, w10, w02, w20, w03, w30;
    wire [7:0] w12, w21, w13, w31, w23, w32;

    recurrent_layer uut (
        .clk(clk), .rst_n(rst_n), .ext_spike_in(ext_in),
        .spike_out(spk),
        .v_mem_0(v0), .v_mem_1(v1), .v_mem_2(v2), .v_mem_3(v3),
        .w01(w01), .w10(w10), .w02(w02), .w20(w20),
        .w03(w03), .w30(w30), .w12(w12), .w21(w21),
        .w13(w13), .w31(w31), .w23(w23), .w32(w32)
    );

    initial clk = 0;
    always #5 clk = ~clk;

    task tick;
        input [3:0] pattern;
        begin
            @(posedge clk); #1;
            ext_in = pattern;
        end
    endtask

    integer i;
    initial begin
        $dumpfile("recurrent_dump.vcd");
        $dumpvars(0, tb_recurrent_layer);

        rst_n  = 0; ext_in = 4'b0000;
        @(posedge clk); #1;
        @(posedge clk); #1;
        rst_n = 1;

        // =====================================================================
        // [Phase 1] 베이스라인: N0만 자극 → N0만 발화하는지 확인
        // =====================================================================
        $display("\n=== [Phase 1] 베이스라인: N0만 자극 (학습 전) ===");
        $display("기대: N0만 발화, N1은 발화 안 함");
        for (i = 0; i < 10; i = i + 1)
            tick(4'b0001); // N0만 자극
        tick(4'b0000);

        // =====================================================================
        // [Phase 2] 패턴 A 학습: N0+N1 동시 자극 50회
        //   → W01, W10 강화 기대
        // =====================================================================
        $display("\n=== [Phase 2] 패턴 A 학습: N0+N1 동시 자극 50회 ===");
        $display("W01, W10이 5에서 증가하면 학습 성공!");
        for (i = 0; i < 50; i = i + 1)
            tick(4'b0011); // N0+N1 동시 자극
        tick(4'b0000);

        // 안정화 대기
        for (i = 0; i < 10; i = i + 1)
            tick(4'b0000);

        // =====================================================================
        // [Phase 3] 연상 복원: N0만 자극
        //   → 학습된 W01으로 N1도 발화하는지 확인
        //   → 이것이 "연상 기억 (Associative Memory)"
        // =====================================================================
        $display("\n=== [Phase 3] 연상 복원: N0만 자극 (학습 후) ===");
        $display("기대: N0 발화 → W01 강화 → N1도 발화! (패턴 복원)");
        for (i = 0; i < 20; i = i + 1)
            tick(4'b0001); // N0만 자극
        tick(4'b0000);

        // =====================================================================
        // [Phase 4] 패턴 B 학습: N2+N3 동시 자극
        //   → W23, W32 강화 (패턴 A와 독립적)
        // =====================================================================
        $display("\n=== [Phase 4] 패턴 B 학습: N2+N3 동시 자극 ===");
        for (i = 0; i < 50; i = i + 1)
            tick(4'b1100); // N2+N3 동시 자극
        tick(4'b0000);

        for (i = 0; i < 5; i = i + 1)
            tick(4'b0000);

        // =====================================================================
        // [Phase 5] 패턴 B 복원: N2만 자극
        //   → N3도 발화하는지 확인
        // =====================================================================
        $display("\n=== [Phase 5] 패턴 B 복원: N2만 자극 ===");
        $display("기대: N2 발화 → N3도 발화! (패턴 B 복원)");
        for (i = 0; i < 20; i = i + 1)
            tick(4'b0100); // N2만 자극

        $display("\n=== [시뮬레이션 완료] ===");
        $finish;
    end

    // 핵심 시냅스 가중치와 발화 패턴 모니터링
    initial begin
        $monitor("T=%t | In=%b | Spk=%b | V0=%3d V1=%3d V2=%3d V3=%3d | W01=%3d W10=%3d W23=%3d W32=%3d",
                 $time, ext_in, spk, v0, v1, v2, v3, w01, w10, w23, w32);
    end

endmodule
// =============================================================================
// End of tb_recurrent_layer.v
// =============================================================================
