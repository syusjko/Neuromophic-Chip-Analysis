// =============================================================================
// Module  : tb_lif_neuron (Testbench)
// Description : lif_neuron 모듈에 입력을 주어 파형을 관찰하는 시뮬레이션 코드
//
// [수정 사항]
//   1. spike_in 할당을 클럭 엣지 '이전'에 설정 (#1 딜레이 기법 사용)
//      → @(posedge clk) 이후 #1을 주어 셋업 타임 위반 없이 다음 클럭에 반영
//   2. 시나리오 1의 repeat 횟수를 30으로 늘려 확실한 발화 유도
//   3. 발화 후 리셋 동작 확인 시나리오 추가
// =============================================================================
`timescale 1ns / 1ps

module tb_lif_neuron;

    // -------------------------------------------------------------------------
    // 1. 신호 선언
    // -------------------------------------------------------------------------
    reg        clk;
    reg        rst_n;
    reg        spike_in;

    wire       spike_out;
    wire [7:0] v_mem;

    // -------------------------------------------------------------------------
    // 2. DUT (Device Under Test) 연결
    //    THRESHOLD=60으로 낮춰서 빠른 발화 확인
    // -------------------------------------------------------------------------
    lif_neuron #(
        .THRESHOLD(8'd60),
        .LEAK     (8'd5),
        .WEIGHT   (8'd10)
    ) uut (
        .clk      (clk),
        .rst_n    (rst_n),
        .spike_in (spike_in),
        .spike_out(spike_out),
        .v_mem    (v_mem)
    );

    // -------------------------------------------------------------------------
    // 3. 클럭 생성 (10ns 주기 = 100MHz)
    // -------------------------------------------------------------------------
    initial clk = 0;
    always  #5 clk = ~clk;

    // -------------------------------------------------------------------------
    // 4. 태스크 정의: 클럭 엣지 이후 #1 딜레이로 spike_in 안전하게 설정
    //    → 시뮬레이터의 race condition 방지 (Non-blocking 관행)
    // -------------------------------------------------------------------------
    task set_spike;
        input val;
        begin
            @(posedge clk);
            #1;              // 클럭 엣지 직후 1ns 딜레이 → 다음 클럭에 확실히 반영
            spike_in = val;
        end
    endtask

    // -------------------------------------------------------------------------
    // 5. 시뮬레이션 시나리오
    // -------------------------------------------------------------------------
    integer i;

    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, tb_lif_neuron);

        // --- 초기화 ---
        rst_n    = 0;
        spike_in = 0;

        // 리셋 2클럭 유지 후 해제
        @(posedge clk); #1;
        @(posedge clk); #1;
        rst_n = 1;

        // =================================================================
        // [시나리오 1] 연속 스파이크 입력 → 발화(Firing) 유도
        //   THRESHOLD=60, 순증가=WEIGHT-LEAK=5/cycle
        //   → 60/5 = 12 클럭 이상이면 발화 예상
        //   30클럭 연속 입력 → 발화 후 리셋까지 관찰
        // =================================================================
        $display("\n[시나리오 1] 연속 스파이크 30회 입력 (발화 유도)");
        for (i = 0; i < 30; i = i + 1) begin
            set_spike(1);
        end

        // =================================================================
        // [시나리오 2] 입력 중단 → Leak 동작 확인 (전압 선형 감소)
        // =================================================================
        $display("\n[시나리오 2] 입력 중단 → Leak 감소 관찰");
        for (i = 0; i < 10; i = i + 1) begin
            set_spike(0);
        end

        // =================================================================
        // [시나리오 3] 재입력 → 두 번째 발화 확인
        // =================================================================
        $display("\n[시나리오 3] 재입력 → 두 번째 발화 확인");
        for (i = 0; i < 20; i = i + 1) begin
            set_spike(1);
        end

        // =================================================================
        // [시나리오 4] 입력 중단 → Underflow 방지 확인 (0 이하로 안 내려감)
        // =================================================================
        $display("\n[시나리오 4] 입력 중단 → Underflow 방지 확인");
        for (i = 0; i < 20; i = i + 1) begin
            set_spike(0);
        end

        // =================================================================
        // [시나리오 5] 리셋 동작 확인
        // =================================================================
        $display("\n[시나리오 5] 리셋 동작 확인");
        // 전압 어느 정도 올린 뒤
        for (i = 0; i < 5; i = i + 1) begin
            set_spike(1);
        end
        // 리셋 인가
        @(posedge clk); #1;
        rst_n = 0;
        @(posedge clk); #1;
        @(posedge clk); #1;
        rst_n = 1;
        // 리셋 후 전압이 0인지 확인
        for (i = 0; i < 3; i = i + 1) begin
            set_spike(0);
        end

        #20;
        $display("\n[시뮬레이션 완료]");
        $finish;
    end

    // -------------------------------------------------------------------------
    // 6. 모니터링
    // -------------------------------------------------------------------------
    initial begin
        $monitor("Time=%t | Input=%b | Voltage=%3d | Fired?=%b",
                 $time, spike_in, v_mem, spike_out);
    end

endmodule
// =============================================================================
// End of tb_lif_neuron.v
// =============================================================================
