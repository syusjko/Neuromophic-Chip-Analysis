// =============================================================================
// Module  : tb_network (v3 - STDP 학습 버그 수정)
//
// [버그 수정]
//   기존 파라미터 문제:
//     N1 발화 주기 = 5클럭, 그 사이 N2 Leak = -5 × 5 = -25
//     N1 발화 시 N2에 전달되는 전류 = weight(10) → 누적 불가능
//     → N2가 절대 발화 못함 → post_spike=0 → LTP 조건 불성립 → weight 고정
//
//   해결책:
//     N2_LEAK=1로 줄여 전압 유지 시간 연장
//     SYN_INIT_WEIGHT=30으로 올려 N2가 초반에 발화 가능하게
//     → N2 발화 후 LTP 적용 → weight 증가 → 더 빠른 발화 확인
//
// 관전 포인트:
//   Syn_W가 30 → 32 → 34 ... 증가하면 STDP LTP 학습 성공!
//   N2 발화 주기가 점점 짧아지면 완벽!
// =============================================================================
`timescale 1ns / 1ps

module tb_network;

    // -------------------------------------------------------------------------
    // 신호 선언
    // -------------------------------------------------------------------------
    reg        clk;
    reg        rst_n;
    reg        spike_in;

    wire       spike_out_n1;
    wire       spike_out_n2;
    wire [7:0] v1, v2;
    wire [7:0] syn_weight;

    // -------------------------------------------------------------------------
    // DUT 연결 (파라미터 재설계)
    //
    // N1: THRESHOLD=60, LEAK=5, INPUT_CURRENT=20
    //     → 순증가 +15/cycle → 4클럭마다 발화
    //
    // Synapse: INIT_WEIGHT=30
    //     → N1 발화 시 N2에 30 전달
    //
    // N2: THRESHOLD=60, LEAK=1
    //     → N1 발화 사이 4클럭 동안 Leak = -1×4 = -4 (매우 적음)
    //     → 30 → 26 → 22 → 18 → 14 (다음 N1 발화) → 44 → ...
    //     → 2번째 N1 발화 후: 44 → 40 → 36 → 32 → 28 (다음) → 58
    //     → 3번째 N1 발화 후: 58 → 54 → 50 → 46 → 42 (다음) → 72 > 60 → 발화!
    // -------------------------------------------------------------------------
    network #(
        .N1_THRESHOLD    (8'd60),
        .N1_LEAK         (8'd5),
        .N1_INPUT_CURRENT(8'd20),
        .N2_THRESHOLD    (8'd60),
        .N2_LEAK         (8'd1),   // ← 핵심 수정: Leak 줄여서 N2 전압 유지
        .SYN_INIT_WEIGHT (8'd30),  // ← 핵심 수정: 초기 weight 높여서 N2 발화 유도
        .SYN_LTP_STEP    (8'd2),   // LTP 스텝 2 (학습 효과 빠르게 관찰)
        .SYN_LTD_STEP    (8'd1),
        .SYN_TRACE_DECAY (4'd8)
    ) uut (
        .clk            (clk),
        .rst_n          (rst_n),
        .spike_in_global(spike_in),
        .spike_out_n1   (spike_out_n1),
        .spike_out_n2   (spike_out_n2),
        .v_mem_n1       (v1),
        .v_mem_n2       (v2),
        .syn_weight     (syn_weight)
    );

    // -------------------------------------------------------------------------
    // 클럭 생성 (10ns = 100MHz)
    // -------------------------------------------------------------------------
    initial clk = 0;
    always  #5 clk = ~clk;

    // -------------------------------------------------------------------------
    // 태스크
    // -------------------------------------------------------------------------
    task set_spike;
        input val;
        begin
            @(posedge clk); #1;
            spike_in = val;
        end
    endtask

    integer i;

    initial begin
        $dumpfile("network_dump.vcd");
        $dumpvars(0, tb_network);

        rst_n    = 0;
        spike_in = 0;
        @(posedge clk); #1;
        @(posedge clk); #1;
        rst_n = 1;

        // =================================================================
        // [시나리오 1] 연속 자극 150회
        //   초반: weight=30 → N2가 3~4번 N1 발화 후 첫 발화
        //   LTP 적용 후: weight 증가 → N2 발화 주기 단축 확인
        // =================================================================
        $display("\n[시나리오 1] 연속 자극 150회 - STDP LTP 학습 관찰");
        $display("  Syn_W가 30에서 증가하면 학습 성공!");
        for (i = 0; i < 150; i = i + 1) begin
            set_spike(1);
        end

        // =================================================================
        // [시나리오 2] 입력 중단 - Leak 관찰 (weight는 유지됨)
        // =================================================================
        $display("\n[시나리오 2] 입력 중단 - weight 유지 확인");
        for (i = 0; i < 20; i = i + 1) begin
            set_spike(0);
        end

        // =================================================================
        // [시나리오 3] 재자극 - 학습된 weight로 N2 더 빨리 발화하는지 확인
        // =================================================================
        $display("\n[시나리오 3] 재자극 - 높아진 weight 효과 확인");
        for (i = 0; i < 80; i = i + 1) begin
            set_spike(1);
        end

        $display("\n[시뮬레이션 완료]");
        $finish;
    end

    // -------------------------------------------------------------------------
    // 모니터링
    // -------------------------------------------------------------------------
    initial begin
        $monitor("T=%t | In=%b | N1_V=%3d(F:%b) | Syn_W=%3d | N2_V=%3d(F:%b)",
                 $time, spike_in,
                 v1, spike_out_n1,
                 syn_weight,
                 v2, spike_out_n2);
    end

endmodule
// =============================================================================
// End of tb_network.v (v3)
// =============================================================================
